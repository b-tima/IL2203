library verilog;
use verilog.vl_types.all;
entity svtb is
end svtb;
