library IEEE;
use ieee.std_logic_1164.all;

entity test is port(); end test;