library verilog;
use verilog.vl_types.all;
entity svtb_sv_unit is
end svtb_sv_unit;
